
module system (
	clk_clk,
	reset_reset_n,
	parallelport_0_conduit_parport_export);	

	input		clk_clk;
	input		reset_reset_n;
	inout	[7:0]	parallelport_0_conduit_parport_export;
endmodule
