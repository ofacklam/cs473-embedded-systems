
module system (
	clk_clk,
	reset_reset_n,
	customuart_0_trx_out_rx,
	customuart_0_trx_out_tx);	

	input		clk_clk;
	input		reset_reset_n;
	input		customuart_0_trx_out_rx;
	output		customuart_0_trx_out_tx;
endmodule
